magic
tech gf180mcuD
timestamp 1755274543
<< nwell >>
rect -33 -57 150 14
<< nmos >>
rect 12 -102 18 -85
rect 39 -102 45 -85
rect 63 -102 69 -85
rect 92 -102 98 -85
<< pmos >>
rect 12 -43 18 -9
rect 39 -43 45 -9
rect 63 -43 69 -9
rect 92 -43 98 -9
<< ndiff >>
rect -6 -87 12 -85
rect -6 -93 1 -87
rect 8 -93 12 -87
rect -6 -102 12 -93
rect 18 -102 39 -85
rect 45 -102 63 -85
rect 69 -102 92 -85
rect 98 -89 122 -85
rect 98 -95 110 -89
rect 116 -95 122 -89
rect 98 -102 122 -95
<< pdiff >>
rect -4 -14 12 -9
rect -4 -31 -2 -14
rect 8 -31 12 -14
rect -4 -43 12 -31
rect 18 -15 39 -9
rect 18 -32 25 -15
rect 35 -32 39 -15
rect 18 -43 39 -32
rect 45 -11 63 -9
rect 45 -28 49 -11
rect 59 -28 63 -11
rect 45 -43 63 -28
rect 69 -16 92 -9
rect 69 -33 75 -16
rect 85 -33 92 -16
rect 69 -43 92 -33
rect 98 -14 119 -9
rect 98 -31 104 -14
rect 114 -31 119 -14
rect 98 -43 119 -31
<< ndiffc >>
rect 1 -93 8 -87
rect 110 -95 116 -89
<< pdiffc >>
rect -2 -31 8 -14
rect 25 -32 35 -15
rect 49 -28 59 -11
rect 75 -33 85 -16
rect 104 -31 114 -14
<< psubdiff >>
rect -30 -104 -17 -102
rect -30 -111 -28 -104
rect -19 -111 -17 -104
rect 134 -106 148 -104
rect -30 -114 -17 -111
rect 134 -111 137 -106
rect 145 -111 148 -106
rect 134 -113 148 -111
<< nsubdiff >>
rect -4 8 9 11
rect -4 2 -1 8
rect 5 2 9 8
rect 103 7 115 10
rect -4 0 9 2
rect 103 1 106 7
rect 112 1 115 7
rect 103 -1 115 1
<< psubdiffcont >>
rect -28 -111 -19 -104
rect 137 -111 145 -106
<< nsubdiffcont >>
rect -1 2 5 8
rect 106 1 112 7
<< polysilicon >>
rect 12 -9 18 4
rect 39 -9 45 5
rect 63 -9 69 5
rect 92 -9 98 5
rect 12 -57 18 -43
rect 3 -60 18 -57
rect 3 -65 7 -60
rect 15 -65 18 -60
rect 3 -67 18 -65
rect 12 -85 18 -67
rect 39 -69 45 -43
rect 31 -71 45 -69
rect 31 -77 34 -71
rect 41 -77 45 -71
rect 31 -79 45 -77
rect 39 -85 45 -79
rect 63 -58 69 -43
rect 63 -60 76 -58
rect 63 -65 66 -60
rect 74 -65 76 -60
rect 63 -68 76 -65
rect 63 -85 69 -68
rect 92 -73 98 -43
rect 92 -75 107 -73
rect 92 -80 98 -75
rect 104 -80 107 -75
rect 92 -83 107 -80
rect 92 -85 98 -83
rect 12 -107 18 -102
rect 39 -107 45 -102
rect 63 -108 69 -102
rect 92 -107 98 -102
<< polycontact >>
rect 7 -65 15 -60
rect 34 -77 41 -71
rect 66 -65 74 -60
rect 98 -80 104 -75
<< metal1 >>
rect -13 8 120 14
rect -13 2 -1 8
rect 5 7 120 8
rect 5 2 106 7
rect -13 1 106 2
rect 112 1 120 7
rect -13 -1 120 1
rect -3 -14 9 -1
rect 48 -11 60 -1
rect -3 -31 -2 -14
rect 8 -31 9 -14
rect -3 -32 9 -31
rect 24 -15 36 -13
rect 24 -32 25 -15
rect 35 -32 36 -15
rect 48 -28 49 -11
rect 59 -28 60 -11
rect 102 -14 115 -1
rect 48 -30 60 -28
rect 74 -16 86 -15
rect 24 -39 36 -32
rect 74 -33 75 -16
rect 85 -33 86 -16
rect 74 -39 86 -33
rect 102 -31 104 -14
rect 114 -31 115 -14
rect 102 -37 115 -31
rect 24 -43 86 -39
rect 24 -49 49 -43
rect 58 -49 86 -43
rect 24 -53 86 -49
rect 3 -59 18 -57
rect 3 -65 7 -59
rect 15 -65 18 -59
rect 3 -67 18 -65
rect 31 -71 45 -69
rect 31 -77 34 -71
rect 42 -77 45 -71
rect 31 -79 45 -77
rect 50 -86 59 -53
rect 64 -60 76 -58
rect 64 -66 66 -60
rect 74 -66 76 -60
rect 64 -67 76 -66
rect 93 -75 107 -73
rect 93 -81 97 -75
rect 105 -81 107 -75
rect 93 -82 107 -81
rect -1 -87 59 -86
rect -1 -93 1 -87
rect 8 -93 59 -87
rect -1 -94 59 -93
rect 106 -89 119 -87
rect -1 -95 57 -94
rect 106 -95 110 -89
rect 116 -95 119 -89
rect 106 -101 119 -95
rect -32 -104 150 -101
rect -32 -111 -28 -104
rect -19 -106 150 -104
rect -19 -111 137 -106
rect 145 -111 150 -106
rect -32 -116 150 -111
<< via1 >>
rect 49 -49 58 -43
rect 7 -60 15 -59
rect 7 -65 15 -60
rect 34 -77 41 -71
rect 41 -77 42 -71
rect 66 -65 74 -60
rect 66 -66 74 -65
rect 97 -80 98 -75
rect 98 -80 104 -75
rect 104 -80 105 -75
rect 97 -81 105 -80
<< metal2 >>
rect 47 -43 60 -40
rect 47 -49 49 -43
rect 58 -49 60 -43
rect 47 -52 60 -49
rect 6 -59 17 -57
rect 6 -65 7 -59
rect 15 -65 17 -59
rect 6 -66 17 -65
rect 64 -60 76 -58
rect 64 -66 66 -60
rect 74 -66 76 -60
rect 64 -68 76 -66
rect 32 -71 44 -69
rect 32 -77 34 -71
rect 42 -77 44 -71
rect 32 -79 44 -77
rect 93 -75 108 -73
rect 93 -81 97 -75
rect 105 -81 108 -75
rect 93 -82 108 -81
<< labels >>
rlabel metal1 5 -1 106 14 0 VDD
rlabel metal1 -19 -116 137 -101 0 VSS
rlabel metal1 0 0 0 0 0 Y
rlabel polycontact 7 -65 15 -60 0 A
rlabel polysilicon 34 -77 42 -71 0 B
rlabel polycontact 66 -65 74 -60 0 C
rlabel polycontact 98 -80 104 -75 0 D
<< end >>
