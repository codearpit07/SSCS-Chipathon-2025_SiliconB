* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__nand4_1.ext - technology: gf180mcuD

.subckt gf180mcu_osu_sc_gp9t3v3__nand4_1 A B C D Y VDD VSS

X0 Y A VDD VDD pfet_03v3 W=1.70000U L=0.300000U
X1 Y B VDD VDD pfet_03v3 W=1.70000U L=0.300000U
X2 Y C VDD VDD pfet_03v3 W=1.70000U L=0.300000U
X3 Y D VDD VDD pfet_03v3 W=1.70000U L=0.300000U
X4 Y A net1 VSS nfet_03v3 W=0.850000U L=0.300000U
X5 net1 B net2 VSS nfet_03v3 W=0.850000U L=0.300000U
X6 net2 C net3 VSS nfet_03v3 W=0.850000U L=0.300000U
X7 net3 D VSS VSS nfet_03v3 W=0.850000U L=0.300000U

.ends
