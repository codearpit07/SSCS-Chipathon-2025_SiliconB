magic
tech gf180mcuD
timestamp 1755276715
<< nwell >>
rect -6 23 78 75
<< nmos >>
rect 15 -23 21 -6
rect 33 -23 39 -6
rect 51 -23 57 -6
<< pmos >>
rect 15 32 21 66
rect 33 32 39 66
rect 51 32 57 66
<< ndiff >>
rect 3 -11 15 -6
rect 3 -19 6 -11
rect 11 -19 15 -11
rect 3 -23 15 -19
rect 21 -11 33 -6
rect 21 -19 24 -11
rect 29 -19 33 -11
rect 21 -23 33 -19
rect 39 -11 51 -6
rect 39 -19 42 -11
rect 47 -19 51 -11
rect 39 -23 51 -19
rect 57 -11 69 -6
rect 57 -19 60 -11
rect 65 -19 69 -11
rect 57 -23 69 -19
<< pdiff >>
rect 3 56 15 66
rect 3 40 6 56
rect 11 40 15 56
rect 3 32 15 40
rect 21 56 33 66
rect 21 40 24 56
rect 29 40 33 56
rect 21 32 33 40
rect 39 56 51 66
rect 39 40 42 56
rect 47 40 51 56
rect 39 32 51 40
rect 57 56 69 66
rect 57 40 60 56
rect 65 40 69 56
rect 57 32 69 40
<< ndiffc >>
rect 6 -19 11 -11
rect 24 -19 29 -11
rect 42 -19 47 -11
rect 60 -19 65 -11
<< pdiffc >>
rect 6 40 11 56
rect 24 40 29 56
rect 42 40 47 56
rect 60 40 65 56
<< psubdiff >>
rect -4 -32 13 -30
rect -4 -38 0 -32
rect 8 -38 13 -32
rect -4 -42 13 -38
rect 26 -32 43 -30
rect 26 -38 31 -32
rect 39 -38 43 -32
rect 26 -42 43 -38
rect 60 -32 77 -30
rect 60 -38 65 -32
rect 73 -38 77 -32
rect 60 -42 77 -38
<< nsubdiff >>
rect -5 86 12 88
rect -5 80 -2 86
rect 6 80 12 86
rect -5 76 12 80
rect 27 86 44 88
rect 27 80 31 86
rect 39 80 44 86
rect 27 76 44 80
rect 60 86 77 88
rect 60 80 64 86
rect 72 80 77 86
rect 60 76 77 80
<< psubdiffcont >>
rect 0 -38 8 -32
rect 31 -38 39 -32
rect 65 -38 73 -32
<< nsubdiffcont >>
rect -2 80 6 86
rect 31 80 39 86
rect 64 80 72 86
<< polysilicon >>
rect 15 66 21 73
rect 33 66 39 73
rect 51 66 57 73
rect 15 5 21 32
rect 33 21 39 32
rect 30 19 39 21
rect 30 14 32 19
rect 37 14 39 19
rect 30 12 39 14
rect 9 3 21 5
rect 9 -2 11 3
rect 16 -2 21 3
rect 9 -4 21 -2
rect 15 -6 21 -4
rect 33 -6 39 12
rect 51 5 57 32
rect 45 3 57 5
rect 45 -2 47 3
rect 52 -2 57 3
rect 45 -4 57 -2
rect 51 -6 57 -4
rect 15 -28 21 -23
rect 33 -28 39 -23
rect 51 -28 57 -23
<< polycontact >>
rect 32 14 37 19
rect 11 -2 16 3
rect 47 -2 52 3
<< metal1 >>
rect -6 86 78 88
rect -6 80 -2 86
rect 6 80 31 86
rect 39 80 64 86
rect 72 80 78 86
rect -6 72 78 80
rect 5 67 49 72
rect 5 56 13 67
rect 5 40 6 56
rect 11 40 13 56
rect 5 36 13 40
rect 23 56 31 62
rect 23 40 24 56
rect 29 40 31 56
rect 23 31 31 40
rect 41 56 49 67
rect 41 40 42 56
rect 47 40 49 56
rect 41 36 49 40
rect 59 56 67 62
rect 59 40 60 56
rect 65 40 67 56
rect 59 31 67 40
rect 23 29 67 31
rect 23 28 71 29
rect 23 26 63 28
rect 59 22 63 26
rect 70 22 71 28
rect 59 21 71 22
rect 30 20 39 21
rect 30 14 31 20
rect 38 14 39 20
rect 30 12 39 14
rect 9 4 18 5
rect 9 -2 10 4
rect 17 -2 18 4
rect 9 -4 18 -2
rect 45 4 54 5
rect 45 -2 46 4
rect 53 -2 54 4
rect 45 -4 54 -2
rect 5 -11 13 -9
rect 5 -19 6 -11
rect 11 -19 13 -11
rect 5 -26 13 -19
rect 23 -11 31 -9
rect 23 -19 24 -11
rect 29 -19 31 -11
rect 23 -21 31 -19
rect 41 -11 49 -9
rect 41 -19 42 -11
rect 47 -19 49 -11
rect 41 -21 49 -19
rect 59 -11 67 21
rect 59 -19 60 -11
rect 65 -19 67 -11
rect 59 -21 67 -19
rect -6 -32 78 -26
rect -6 -38 0 -32
rect 8 -38 31 -32
rect 39 -38 65 -32
rect 73 -38 78 -32
rect -6 -42 78 -38
<< via1 >>
rect 63 22 70 28
rect 31 19 38 20
rect 31 14 32 19
rect 32 14 37 19
rect 37 14 38 19
rect 10 3 17 4
rect 10 -2 11 3
rect 11 -2 16 3
rect 16 -2 17 3
rect 46 3 53 4
rect 46 -2 47 3
rect 47 -2 52 3
rect 52 -2 53 3
<< metal2 >>
rect 62 28 71 29
rect 62 22 63 28
rect 70 22 71 28
rect 62 21 71 22
rect 30 20 39 21
rect 30 14 31 20
rect 38 14 39 20
rect 30 12 39 14
rect 9 4 18 5
rect 9 -2 10 4
rect 17 -2 18 4
rect 9 -4 18 -2
rect 45 4 54 5
rect 45 -2 46 4
rect 53 -2 54 4
rect 45 -4 54 -2
<< labels >>
rlabel metal2 51 1 52 2 1 A
rlabel metal2 34 17 35 18 1 B
rlabel metal2 14 1 15 2 1 C
rlabel via1 66 26 67 27 1 Y
<< end >>
